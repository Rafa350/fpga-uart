module UART_RX
(
    input  logic       i_clock,
    input  logic       i_reset,

    output logic [7:0] o_data);

endmodule